magic
tech scmos
timestamp 1596723265
<< nwell >>
rect -4 3 17 24
<< polysilicon >>
rect 3 11 7 13
rect 3 -2 7 6
rect 2 -6 7 -2
rect 3 -8 7 -6
rect 3 -20 7 -18
<< ndiffusion >>
rect -4 -13 3 -8
rect -4 -18 -2 -13
rect 2 -18 3 -13
rect 7 -13 8 -8
rect 7 -18 12 -13
<< pdiffusion >>
rect 2 6 3 11
rect 7 6 8 11
<< metal1 >>
rect -2 22 15 23
rect -2 17 -1 22
rect 4 17 9 22
rect 14 17 15 22
rect -2 15 15 17
rect -2 11 2 15
rect 8 1 12 6
rect -7 -2 0 -1
rect -7 -6 -3 -2
rect 8 -4 24 1
rect -7 -7 0 -6
rect 8 -8 12 -4
rect -2 -21 2 -18
rect -2 -22 15 -21
rect -2 -27 -1 -22
rect 4 -27 9 -22
rect 14 -27 15 -22
rect -2 -28 15 -27
<< ntransistor >>
rect 3 -18 7 -8
<< ptransistor >>
rect 3 6 7 11
<< polycontact >>
rect -3 -6 2 -2
<< ndcontact >>
rect -2 -18 2 -13
rect 8 -13 12 -8
<< pdcontact >>
rect -2 6 2 11
rect 8 6 12 11
<< psubstratepcontact >>
rect -1 -27 4 -22
rect 9 -27 14 -22
<< nsubstratencontact >>
rect -1 17 4 22
rect 9 17 14 22
<< labels >>
rlabel metal1 -2 23 15 23 5 VDD
rlabel metal1 -2 -28 15 -28 1 Ground
rlabel metal1 23 -4 23 1 7 Vout
rlabel metal1 -6 -7 -6 -1 3 Vin
<< end >>
